/*
This system verilog module performs the functionality of instruction decoder
Author : Anindya Kishore Choudhury (anindyakchoudhury@gmail.com)
*/

`include "simple_processor_pkg.sv"

module ins_dec
import simple_processor_pkg::*;
#(
    //-PARAMETERS
    //-LOCALPARAMS
) (
    //-PORTS
    input  logic [INSTR_WIDTH-1:0] imem_rdata_i, //instruction data coming from IMEM
    input  logic                   imem_ack_i,   //IMEM acknowledge to select between imem_rdata_i or 0

    output func_t                  func_o,       //op codes are stored in this typedef
    output logic                   we_o,         //write enable pin
    output logic [2:0]             rd_addr_o,    //destination register address
    output logic [2:0]             rs1_addr_o,   //RS1 register address
    output logic [2:0]             rs2_addr_o,   //RS2 register address
    output logic [5:0]             imm_o,        //unextended immediate
    output logic                   valid_pc      //for mux selector input after pc
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic [INSTR_WIDTH-1:0] instruction;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign instruction = imem_ack_i ? imem_rdata_i : '0;
  assign func_o      = instruction[3:0];
  assign rs1_addr_o  = instruction[12:10];
  assign imm_o       = instruction[9:4];
  assign rs2_addr_o  = instruction[9:7];
  assign rd_addr_o   = instruction[15:13]

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (DATA_WIDTH > 2) begin
      $display("\033[1;33m%m DATA_WIDTH\033[0m");
    end
  end
`endif  // SIMULATION

endmodule
