git /*
Write a markdown documentation for this systemverilog module:
Author :  ()
*/

module FIFO_ANJAN #(
    Data_width=8
    Mem_Depth=16
//-PARAMETERS
    //-LOCALPARAMS
) (
input logic clk_i,
input logic arst_ni,
input logic ,boot_addr_i,
output logic imem_req_odmem_ack_i, 
output logic imem_addr_o,
output logic dmem_req_o,
output logic dmem_wr_o,
output logic dmem_addr_o,
output logic dmem_wdata_o,
output logic ddmem_rdata_i,
output logic dmem_ack_i,
input logic  imem_rdata_i,
input logic imem_ack_i ,
//-PORTS
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////
 logic [FIFO_SIZE:0] wr_ptr;
 logic [FIFO_SIZE:0] rd_ptr;
 logic [FIFO_SIZE:0] wr_ptr_next;
 logic [FIFO_SIZE:0] rd_ptr_next;
 logic hsi;
 logic hso;
 logic msb_eq;
 logic nmsb_eq;
 logic empty;
 logic full;

 logic [ELEM_WIDTH-1:0] elem_out;
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////
 assign hsi=elem_in_valid_i & elem_in_ready_o;
 assign hso=elem_out_valid_o & elem_out_ready_i;

 always_ff @(posedge clk or negedge rstn)
  
 if (hsi && rd_ptr<=3)
  rd_ptr=rd_ptr+1;
  else
    rd_ptr=0;
  if (hso &&)
    wr_ptr=wr_ptr+1;
    if 
 
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (DATA_WIDTH > 2) begin
      $display("\033[1;33m%m DATA_WIDTH\033[0m");
    end
  end
`endif  // SIMULATION

endmodule
