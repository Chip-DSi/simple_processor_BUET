/*
Write a markdown documentation for this systemverilog module:
Author : Md. Nayem Hasan (nayem90375@gmail.com)
*/

module alumem
import simple_processor_pkg::DATA_WIDTH;
import simple_processor_pkg::ADDR_WIDTH;
 #(
    //parameter int MEM_ADDR_WIDTH =32,
    //parameter int MEM_DATA_WIDTH =32
    //-LOCALPARAMS
) (
   ////////////////////////
    input logic [DATA_WIDTH-1:0] rs1_data_i,   // Data to be stored (for STORE operation)
    input func_t func_i,                        // Function code to select LOAD or STORE
    input logic [DATA_WIDTH-1:0] rs2_data_i,   // Memory address
    input logic we_i,                          // Write enable signal for memory
    input logic [DATA_WIDTH-1:0] mem_data_i,   // Data read from memory (for LOAD operation)
    output logic [DATA_WIDTH-1:0] result,      // Result (data read from memory for LOAD)
    output logic [DATA_WIDTH-1:0] mem_addr_o,  // Memory address output (for LOAD/STORE)
    output logic [DATA_WIDTH-1:0] mem_data_o,  // Data to be written to memory (for STORE)
    output logic mem_write_o                   // Memory write signal (for STORE)


);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  // Memory control signals
// Memory address and data assignments
    assign mem_addr_o = rs2_data_i;
    assign mem_data_o = rs1_data_i;
    assign rs1_data_i =mem_data_i;

  //////////////////////////////////////////////////////////////////////////////////////////////////
// first mux

// LOAD instruction

// STORE instruction


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  // Mimicking the input mux operation
  // Control logic for LOAD and STORE operations
    always_comb begin
    //mem_write_o = 1'b0;  // normally no memory write operation
      case(func_i)
        LOAD: begin
          result = mem_data_i; // Data read from memory
        end
        STORE: always @(posedge clk_i) begin
         // mem_write_o = we_i;   // Enable memory write based on we_i
          result = mem_data_i;  // Data to be stored to memory
        end
        default: begin
          result = 32'b0; // Default result if no valid operation
        end
      endcase
    end
  endmodule
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
initial begin
  if (DATA_WIDTH > 2) begin
    $display("\033[1;33m%m DATA_WIDTH\033[0m");
  end
end
`endif  // SIMULATION

endmodule



