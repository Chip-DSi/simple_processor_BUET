/*
Description
Author : Mymuna Khatun Sadia (maimuna14400@gmail.com)
*/

module AluGateTestbench_tb;

  `define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"
  `include "simple_processor_pkg.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////
parameter int DATA_WIDTH = 32;
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////
logic [DATA_WIDTH-1:0] rd_data_o;
logic [DATA_WIDTH-1:0] rs1_data_i;
logic [DATA_WIDTH-1:0] rs2_data_i;
logic [DATA_WIDTH-1:0] result;
instr_t                func_o;
  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 5ns, 5ns)

logic                  arst_ni = '1;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
// Instantiate rtl_model
  rtl_model #(
    .DATA_WIDTH(DATA_WIDTH)
) dut (
    .rd_data_i(rd_data_o),
    .rs1_data_i(rs1_data_i),
    .rs2_data_i(rs2_data_i),
    .func_o(func_o)
);


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100ns;
    arst_ni <= 0;
    #100ns;
    arst_ni <= 1;
    #100ns;
  endtask


  
// Initial stimulus
initial begin
  // Test case 1: AND operation
  rs1_data_i <= $urandom;
  rs2_data_i <= $urandom;
  func_o = AND;
  result = rs1_data_i & rs2_data_i;
  #10; // Allow some time for the result to propagate
  check_result("Test Case 1", result);

  // Test case 2: OR operation
  rs1_data_i = $urandom;
  rs2_data_i = $urandom;
  func_o = OR;
  result = rs1_data_i | rs2_data_i;
  #10; // Allow some time for the result to propagate
  check_result("Test Case 2", result);

  // Test case 3: XOR operation
  rs1_data_i = $urandom;
  rs2_data_i = $urandom;
  func_o = XOR;
  result = rs1_data_i ^ rs2_data_i;
  #10; // Allow some time for the result to propagate
  check_result("Test Case 3", result);

  // Test case 4: NOT operation
  rs1_data_i = $urandom;
  rs2_data_i = $urandom;
  func_o = NOT;
  result = rs1_data_i ^ rs2_data_i;
  #10; // Allow some time for the result to propagate
  check_result("Test Case 4", result);
end

// Function to check result and display
function void check_result(string name, logic [DATA_WIDTH-1:0] expected);
  if (rd_data_o === expected) begin
      $display("%s: Passed", name);
  end else begin
      $display("%s: Failed. Expected: %h, Got: %h", name, expected, rd_data_i);
  end
endfunction

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    apply_reset();
    start_clk_i();

    @(posedge clk_i);
    result_print(1, "This is a PASS");
    @(posedge clk_i);
    result_print(0, "And this is a FAIL");

    $finish;

  end

endmodule
