/*
Description
Author : B.M.Emroj Hossain Towfik (towfikemroj701@gmail.com)
*/
include "simple_processor_pkg.sv"
`timescale 1ns / 1ps
module alumemtb;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"
import simple_processor_pkg::*;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

    // Parameters and signals for testbench
    localparam DATA_WIDTH = 32;
    localparam ADDR_WIDTH = 32;

    // Clock signal
    reg clk_i = 0;
    always #5 clk_i = ~clk_i; // Toggle every 5 time units

    // Signals for communication with DUT
    logic [DATA_WIDTH-1:0] rs1_data_i;
    logic func_i;
    logic [DATA_WIDTH-1:0] rs2_data_i;
    logic we_i;
    logic [DATA_WIDTH-1:0] mem_data_i;
    logic [DATA_WIDTH-1:0] result;
    logic [DATA_WIDTH-1:0] mem_addr_o;
    logic [DATA_WIDTH-1:0] mem_data_o;
    logic mem_write_o;

    // Instantiate the module under test (alumem)
    alumem #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH)
    ) dut (
        .rs1_data_i(rs1_data_i),
        .func_i(func_i),
        .rs2_data_i(rs2_data_i),
        .we_i(we_i),
        .mem_data_i(mem_data_i),
        .result(result),
        .mem_addr_o(mem_addr_o),
        .mem_data_o(mem_data_o),
        .mem_write_o(mem_write_o)
    );

    // Random number generator for test vectors
   // randbit rand_gen = new();
    //rand_gen.srandom(time);

    // Testbench initialization
    initial begin
        // Apply random test vectors
        repeat (20) begin // Run for 20 transactions
            // Generate random values for test vectors
            rs1_data_i = $urandom_range(0, $urandom_range(0, (2**DATA_WIDTH)-1));
            func_i = $urandom % 2 ? 1'b1 : 1'b0; // Randomly choose LOAD or STORE operation
            rs2_data_i = $urandom_range(0, (2**ADDR_WIDTH)-1);
            we_i = func_i ? 1'b1 : 1'b0; // Set we_i based on func_i for STORE operation
            mem_data_i = $urandom_range(0, (2**DATA_WIDTH)-1);

            // Display inputs for debug
            $display("Time=%0t - Applying transaction", $time);
            $display("rs1_data_i=%h, func_i=%b, rs2_data_i=%h, we_i=%b, mem_data_i=%h", rs1_data_i, func_i, rs2_data_i, we_i, mem_data_i);

            // Wait for a few cycles before applying next transaction
            #10;
        end

        // End simulation
        $display("Simulation finished.");
        $finish;
    end

    // Monitor for debugging (optional)
    always @(posedge clk_i) begin
        // Display signals of interest on positive edge of clock
        $display("Time=%0t - result=%h, mem_addr_o=%h, mem_data_o=%h, mem_write_o=%b", $time, result, mem_addr_o, mem_data_o, mem_write_o);
    end

endmodule
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
 /* `CREATE_CLK(clk_i, 4ns, 6ns)

  logic arst_ni = 1;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100ns;
    arst_ni <= 0;
    #100ns;
    arst_ni <= 1;
    #100ns;
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    apply_reset();
    start_clk_i();

    @(posedge clk_i);
    result_print(1, "This is a PASS");
    @(posedge clk_i);
    result_print(0, "And this is a FAIL");

    $finish;

  end

endmodule
