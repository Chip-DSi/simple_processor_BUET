/*
Write a markdown documentation for this systemverilog module:
Author : Anindya Kishore Choudhury (anindyakchoudhury@gmail.com)
*/

module anindya_FIFO #(
    parameter bit PIPELINED = 1, //determines whether the fifo is pipelined or not
    parameter int DATA_WIDTH = 8,
    parameter int FIFO_SIZE = 4 //means memory depth
    //-LOCALPARAMS
) (
    input logic clk_i, //inp clock signal
    input logic arst_ni, //async active low reset signal
    //input element
    input logic [DATA_WIDTH-1:0] elem_in_i, 
    input logic                  elem_in_valid_i, //input valid signal
    output logic                 elem_in_ready_o, //input ready signal to indicate FIFO is ready to accept the value or not 
    output logic                 elem_out_valid_o, //input valid signal, indicates whether the input element is valid or not
    input logic                  elem_out_ready_i, //output ready signal, whether FIFO is ready to give the output or not
    output logic [DATA_WIDTH-1:0] elem_out_o, //output element

);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  logic [FIFO_SIZE:0] wr_ptr; //write pointer
  logic [FIFO_SIZE:0] rd_ptr; //read pointer

  logic [FIFO_SIZE:0] wr_ptr_next; //write pointer
  logic [FIFO_SIZE:0] rd_ptr_nxt;

  logic hsi; //input handshake
  logic hso; //output handshake 
  
  logic msb_eq;
  logic nmsb_eq;
  
  logic empty;
  logic full;

  logic [DATA_WIDTH] elem_out;
  

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  
  assign hsi = elem_in_valid_i & elem_in_ready_o;
  assign hso = elem_out_valid_o & elem_out_ready_i;

  assign wr_ptr_next = wr_ptr + 1;
  assign rd_ptr_nxt =  rd_ptr + 1;

  assign msb_eq = (wr_ptr[FIFO_SIZE] == rd_ptr[FIFO_SIZE]);
  assign nmsb_eq = (wr_ptr[FIFO_SIZE-1:0] == rd_ptr[FIFO_size-1:0]);

  assign empty = msb_eq & nmsb_eq;
  assign full = !msb_eq & nmsb_eq;

  assign elem_in_ready_o = full ? elem_out_ready_i : '1;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  
  




  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (DATA_WIDTH > 2) begin
      $display("\033[1;33m%m DATA_WIDTH\033[0m");
    end
  end
`endif  // SIMULATION

endmodule
