/*
Description
Author : MD. Toky Tazwar (toky.tech01t@gmail.com)
*/

`include "simple_processor_pkg.sv"

module alu_math_tb;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  import simple_processor_pkg::*;
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 4ns, 6ns)

  logic arst_ni = 1;

  logic  [DATA_WIDTH-1:0] rs1_data_i;
  func_t                  func_i; //added func_t here by akc
  logic  [5:0]            imm;
  logic  [DATA_WIDTH-1:0] rs2_data_i;
  logic  [DATA_WIDTH-1:0] result;
  logic  [DATA_WIDTH-1:0] temp;
  logic  [DATA_WIDTH-1:0] imm_ext;


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////
  int                    pass;
  int                    fail;

//logic [DATA_WIDTH-1:0] ref_mem        [logic [ADDR_WIDTH-1:0]];
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  alu_math dut ( //wrong name put here before
    .rs1_data_i,
    .func_i,
    .imm,
    .rs2_data_i,
    .result
  );
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  task static start_rand_dvr();
  fork
    forever begin
      rs1_data_i   <= $urandom;
      rs2_data_i  <= $urandom;
      imm  <= $urandom;
      randcase
        5: func_i <= ADDI;
        5: func_i <= ADD;
        5: func_i <= SUB;
       // 1: func_i <= INVALID;
    endcase

      @(posedge clk_i);
    end
  join_none
endtask
assign imm_ext = {{26{imm[5]}}, imm};
// monitor and check
task static start_checking();
  fork
    forever begin
      @(posedge clk_i);
      case(func_i)
      ADDI: temp = imm_ext;
      ADD : temp = rs2_data_i;
      SUB : temp = ~rs2_data_i + 1;
      //every other input selection for different block will be done here
       endcase
      if (result === (rs1_data_i + temp)) pass++;
      else begin
        fail++;
      end
    end
  join_none
endtask

//////////////////////////////////////////////////////////////////////////////////////////////////
//-PROCEDURALS
//////////////////////////////////////////////////////////////////////////////////////////////////


  initial begin  // main initial

    //apply_reset();
    //start_clk_i();
    start_checking();
    start_rand_dvr();

    @(posedge clk_i);
    result_print(1, "This is a PASS");
    @(posedge clk_i);
    result_print(0, "And this is a FAIL");

    $finish;

  end

endmodule