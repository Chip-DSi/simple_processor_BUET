/*
Write a markdown documentation for this systemverilog module:
Author : Bokhtiar Foysol Himon (bokhtiarfoysol@gmail.com)
*/

module shift_left (
    input  logic        clk,
    input  logic [31:0] data_in,
    input  logic [4:0]  shift_amount,  // assuming 5-bit shift amount to cover shift ranges from 0 to 31
    output logic [31:0] data_out
);

    always_ff @(posedge clk) begin
        data_out <= data_in << shift_amount;
    end

endmodule

module alu_shift #(
    //-PARAMETERS
    //-LOCALPARAMS
    parameter int DATA_WIDTH = 32
) (
    //-PORTS
    input logic clk,
    input logic [DATA_WIDTH - 1:0] rs1_i,
    input logic [DATA_WIDTH - 1:0] rs2_i,
    input logic [DATA_WIDTH - 1:0] imm,
    input logic use_imm,
    input logic shift_l

    output logic [DATA_WIDTH - 1:0] rd_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

logic [DATA_WIDTH - 1:0] shift_amount;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////
always_comb begin
    if(use_imm)
        shift_amount = imm;
    else
        shift_amount = rs2_i;
end

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

always_ff @(posedge clk) begin
    if(shift_l)
        rd_o <= rs1_i << shift_amount;
    else
        rd_o <= rs1_i >> shift_amount;
end

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (DATA_WIDTH > 2) begin
      $display("\033[1;33m%m DATA_WIDTH\033[0m");
    end
  end
`endif  // SIMULATION

endmodule