/*
Description
Author : Md. Julkar Naim Joy (naimjoy567@gmail.com)
*/
`include "simple_processor_pkg.sv"
module alu_shift_tb;


//module alu_math_tb;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  import simple_processor_pkg::ADDR_WIDTH;
  import simple_processor_pkg::DATA_WIDTH;
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 4ns, 6ns)

  logic arst_ni = 1;

  logic  [DATA_WIDTH-1:0] rs1_data_i;
  logic  [3:0]            func_i;
  logic  [5:0]            imm;
  logic  [DATA_WIDTH-1:0] rs2_data_i;
  logic  [DATA_WIDTH-1:0] result;
  logic  [DATA_WIDTH-1:0] temp;
  logic                   s_r;


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////
  int                    pass;
  int                    fail;

//logic [DATA_WIDTH-1:0] ref_mem        [logic [ADDR_WIDTH-1:0]];
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  alu_shift_tb mem (
    .rs1_data_i,
    .func_i,
    .imm,
    .rs2_data_i,
    .result
  );
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  task static start_rand_dvr();
  fork
    forever begin
      rs1_data_i   <= $urandom;
      rs2_data_i  <= $urandom;
      imm  <= $urandom & 'h11f;
      rand case
        4: func_i <= SLL;
        4: func_i <= SLLI;
        4: func_i <= SLR;
        4: func_i <= SLRI;
    endcase

      @(posedge clk_i);
    end
  join_none
endtask
assign imm = {{26{imm[5]}}, imm};
// monitor and check
task static start_checking();
  fork
    forever begin
      @(posedge clk_i);
      case(func_i)
        SLLI: temp = imm,
              s_r = '0;
        SLRI: temp = imm,
              s_r = '1;
        SLL : temp = rs2_data_i,
              s_r = '0 ;
        SLR : temp = rs2_data_i,
              s_r = '1;
        //every other input selection for different block will be done here
      endcase
      if(s_r=='1)
        if (result === (rs1_data_i >> temp)) pass++;
        else fail++;
      else begin
        if (result === (rs1_data_i << temp)) pass++;
        else fail++;
      end
    end
  join_none
endtask

//////////////////////////////////////////////////////////////////////////////////////////////////
//-PROCEDURALS
//////////////////////////////////////////////////////////////////////////////////////////////////

initial begin  // main initial

  apply_reset();
  start_clk_i();
  //task static start_checking();
  //task static start_rand_dvr();

  start_checking();
  start_rand_dvr();

  @(posedge clk_i);
  result_print(1, "This is a PASS");
  @(posedge clk_i);
  result_print(0, "And this is a FAIL");

  $finish;

end

endmodule