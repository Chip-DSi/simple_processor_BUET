/*
Description
Author : Anindya Kishore Choudhury (anindyakchoudhury@gmail.com)
*/

module demux_tb;

  `define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int NumElem = 6;
  localparam int ElemWidth = 8;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 4ns, 6ns)

  logic arst_ni = 1;
  logic [$clog2(NumElem)-1:0] s_i;
  logic [ElemWidth-1:0] i_i;
  logic [NumElem-1:0][ElemWidth-1:0] o_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  int pass;
  int fail;

  logic [NumElem-1:0][ElemWidth-1:0] ref_out;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  demux #(
    .NUM_ELEM(NumElem),
    .ELEM_WIDTH(ElemWidth)
  ) u_demux (
    .s_i(s_i),
    .i_i(i_i),
    .o_o(o_o)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100ns;
    arst_ni <= 0;
    #100ns;
    arst_ni <= 1;
    #100ns;
  endtask

    // generate random transactions
  task static start_rand_dvr();
    fork
      forever begin
        s_i <= $urandom_range(0, NumElem-1);
        i_i <= $urandom;
        @(posedge clk_i);
      end
    join_none
  endtask

    // monitor and check
  task static start_checking();
    fork
      forever begin
        @(posedge clk_i);
        ref_out      = '0; //understand the importance of this line
        ref_out[s_i] = i_i;

        if (o_o === ref_out) begin
          pass++;
        end else begin
          fail++;
          $display("Error at time %0t: s_i = %0d, i_i = %0h", $time, s_i, i_i);
          $display("Expected o_o = %0h", ref_out);
          $display("Actual o_o   = %0h", o_o);
        end
      end
    join_none
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    apply_reset();
    start_clk_i();
    @(posedge clk_i);
    // Start random driver and checker
    start_rand_dvr();
    start_checking();

    // Run simulation for 1000 cycles
    repeat (1000)@(posedge clk_i);

    // Print results
    result_print(!fail, $sformatf("demux data flow %0d/%0d", pass, pass + fail));

    $finish;

  end

endmodule
