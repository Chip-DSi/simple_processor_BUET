/*
Description
Author : Anindya Kishore Choudhury (anindyakchoudhury@gmail.com)
*/

module register_tb;

  `define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int ElemWidth = 32;
  localparam bit [ElemWidth-1:0] ResetValue = '0;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 4ns, 6ns)

  logic                        arst_ni = '1;
  logic                        en_i = '0;
  logic [ElemWidth-1:0]       d_i = '0;
  logic [ElemWidth-1:0]       q_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  int                          pass;
  int                          fail;
  logic [ElemWidth-1:0]       ref_data;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  register #(
    .ELEM_WIDTH  (ElemWidth),
    .RESET_VALUE (ResetValue)
) u_register (
    .clk_i,
    .arst_ni,
    .en_i,
    .d_i,
    .q_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
  #100ns;
  arst_ni <= 0;
  ref_data <= ResetValue;
  #100ns;
  arst_ni <= 1;
  #100ns;
  endtask

  // generate random transactions
  task static start_rand_dvr();
    fork
      forever begin
        en_i <= $urandom_range(0, 1);
        d_i <= $urandom;
        @(posedge clk_i);
      end
    join_none
  endtask

  // monitor and check
  task static start_checking();
    fork
      forever begin
        @(posedge clk_i);
        if (q_o === ref_data) begin
          pass++;
        end else begin
          fail++;
          //$display("ERROR: Expected q_o = %h, Got q_o = %h at time %t", expected_q, q_o, $time);
        end

        if (~arst_ni) begin
          ref_data = ResetValue;
        end else if (en_i) begin
          ref_data <= d_i;
        end
      end
    join_none
  endtask
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    apply_reset();
    start_clk_i();

    @(posedge clk_i);

    // Data flow checking
    start_rand_dvr();
    start_checking();
    repeat (1000) @(posedge clk_i);
    result_print(!fail, $sformatf("data flow %0d/%0d", pass, pass + fail));

    $finish;

  end

endmodule
