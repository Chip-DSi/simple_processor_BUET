/*
Write a markdown documentation for this systemverilog module:
Author : Bokhtiar Foysol Himon (bokhtiarfoysol@gmail.com)
*/

module himon_FIFO #(
    //-PARAMETERS
    //-LOCALPARAMS
  parameter int Data_Width = 8,
  parameter int Mem_Depth = 16
) (
    //-PORTS
  input logic clk_i,// clk input
  input logic arst_ni, //asynchronous reset negedge
  input logic [Data_Width-1:0] elem_in_i, //input element
  input logic elem_in_valid_i, //indicates if data is valid
  output logic elem_in_ready_o, //indicates if data is ready

  input logic elem_out_ready_i, 
  output logic elem_out_valid_o,
  output logic [Data_Width-1:0] elem_out_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic [Mem_Depth: 0] wr_ptr;
  logic [Mem_Depth: 0] rd_ptr;


  logic [Mem_Depth: 0] wr_next;
  logic [Mem_Depth: 0] rd_next;

  logic hsin;
  logic hsout;

  logic empty;
  logic full;


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////
 
  assign hsin = elem_in_valid_i & elem_in_ready_o;
  assign hsout = elem_out_valid_o & elem_out_ready_i;

  assign wr_next = wr_ptr + 1;
  assign rd_next = rd_ptr + 1;

  if (wr_ptr[Mem_Depth:0] == rd_ptr[Mem_Depth:0])
    assign empty = 1;
  if ((wr_ptr[Mem_Depth - 2 : 0] == rd_ptr[Mem_Depth - 2 : 0])
    && (wr_ptr[Mem_Depth - 1] != rd_ptr[Mem_Depth - 1]))
    assign full = 1;

  if (full==1)
    assign elem_in_ready_o = elem_out_ready_i;
  else
    assign elem_in_ready_o = '1;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (DATA_WIDTH > 2) begin
      $display("\033[1;33m%m DATA_WIDTH\033[0m");
    end
  end
`endif  // SIMULATION

endmodule
