/*
Write a markdown documentation for this systemverilog module:
Author : name (email)
*/

`include "simple_processor_pkg.sv"
module AluGate
import simple_processor_pkg::DATA_WIDTH;
import simple_processor_pkg::INT_REG_WIDTH;
#(

) (
    //-PORTS
output  logic [DATA_WIDTH-1:0] rd_data_o,
input   logic [DATA_WIDTH-1:0] rs1_data_i,
input   logic [DATA_WIDTH-1:0] rs2_data_i,
input   logic                  func_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////
logic [DATA_WIDTH-1:0] result;
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////
//assign imm_ext = {26'b0, imm_o>>4};

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
always_comb begin
    case (func_o)
      AND:      result = rs1_data_i & rs2_data_i;  // AND operation
      OR:       result = rs1_data_i | rs2_data_i;  // OR operation
      XOR:      result = rs1_data_i ^ rs2_data_i;  // XOR operation
      NOT:      result = ~rs1_data_i;              // NOT operation (only uses rs1_data_i)
      default:  result = {DATA_WIDTH{1'b0}};    // Default case to handle invalid opcodes
    endcase
  end

  // Assign the result to the output port
  assign rd_data_o = result;
  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (INT_REG_WIDTH > 32) begin
      $display("\033[1;33m%m TOO MANY REGISTERS\033[0m");
    end
  end
`endif  // SIMULATION

endmodule
